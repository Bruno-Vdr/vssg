module structures

import os
import time
import term
import constants as cst
import util

/**
 * Blog contains arbitrary topic (subject/category/sub-section). This structure store the list of topics,
 * with title (shown) and creation date (time since epoq).
 */
pub struct TopicItem {
pub mut:
	title  string
	date   i64
	locked bool
}

pub struct Blog {
pub:
	name string
mut:
	topics []TopicItem
}

// Static method to build empty Blog struct
pub fn Blog.new(name string) Blog {
	return Blog{name, []TopicItem{}}
}

// Static method, loading blog file from current directory.
pub fn Blog.load() !Blog {
	if util.where_am_i() != .blog_dir {
		return error('Unable to load ${cst.blog_file}.\n[Hint: Are you in the Blog root\'s directory ?]')
	}

	mut ret := util.load_transform_text_file(cst.blog_file, util.del_empty_and_comments)!
	return parse_blog(ret)
}

// exists check for an existing topic with same title as given. Returns boolean accordingly.
pub fn (b Blog) exists(title string) bool {
	for item in b.topics {
		if item.title == title {
			return true
		}
	}
	return false
}

// delete check for an existing topic with same title as given. Returns boolean accordingly.
pub fn (mut b Blog) delete(title string) ! {
	for index, item in b.topics {
		if item.title == title {
			b.topics.delete(index)
			return
		}
	}
	return error('Topic named "${title}" was not found.')
}

// lock_topic check for an existing topic with same title as given. Returns boolean accordingly.
pub fn (mut b Blog) lock_topic(title string) ! {
	for _, mut item in b.topics {
		if item.title == title {
			item.locked = true
			return
		}
	}
	return error('Topic named "${title}" was not found.')
}

// rename the topic with title by new title. Return error if not found.
pub fn (mut b Blog) rename(title string, new_title string) ! {
	mut found := false
	for mut topic in b.topics {
		if title != topic.title {
			continue
		}
		topic.title = new_title
		found = true
		break
	}
	if !found {
		return error('Topic with title "${title}" was not found.')
	}
}

// get_topics_number return numer of topic inside the blog
pub fn (b Blog) get_topics_number() int {
	return b.topics.len
}

pub fn (mut b Blog) add_topic(name string) {
	b.topics << TopicItem{name, (time.ticks() / 1000) + time.offset(), false}
}

pub fn (b Blog) get_topic(i int) ?TopicItem {
	if i < b.topics.len {
		return b.topics[i]
	}
	return none
}

// Save the blog_file configuration.
pub fn (b Blog) save() ! {
	println('Updating ${cst.blog_file}  file in ' + term.blue('${b.name}'))
	mut file := os.open_file('${cst.blog_file}', 'w+', cst.file_access) or {
		return error('Unable to update ${cst.blog_file}: ${err}. ${@FILE_LINE}')
	}

	defer {
		file.close()
	}

	emit_header(mut file, b)!
	emit_topics(mut file, b)!
}

// emit_header write comments and  header only (no topics) int blog_file.
fn emit_header(mut file os.File, b &Blog) ! {
	date_time := time.now().str()
	file.writeln('#\n# Warning: do not edit this file ! It is dynamically generated by vssg.\n# Created on ${date_time} \n# This file contains blog specific parameters for "${b.name}".\n#') or {
		return error('Unable to write ${cst.blog_file}: ${err}. ${@FILE_LINE}')
	}

	file.writeln('name="${b.name}"') or {
		return error('Unable to write name in ${cst.blog_file}: ${err}. ${@FILE_LINE}')
	}
}

// emit_topics writes topics only into blog_file.
fn emit_topics(mut file os.File, b &Blog) ! {
	// Now list the defined topics
	for t in b.topics {
		file.writeln(
			'topic="${t.title}" [${t.date}] [Locked=${t.locked}] # In directory ./${b.name}/' +
			util.obfuscate(t.title)) or {
			return error('Unable to write ${cst.blog_file}: ${err}. ${@FILE_LINE}')
		}
	}
}

/**
 *  Create the initial blog file, containing only the name. At this time, no topics
 * have been added.
 * Note: This method is called in Init command, from outside the blog directory
 * so the configuration file is created with blog directory prepending. Other
 * commands are run from within the blog root's directory (to differentiate them) and
 * access to config_file don't need root's blog prefix.
 */
pub fn (b Blog) create() ! {
	println('Creating ${cst.blog_file}  file in ' + term.blue('${b.name}'))
	mut file := os.open_file('${b.name}${os.path_separator}${cst.blog_file}', 'w+', cst.file_access) or {
		return error('Unable to update ${b.name}${os.path_separator}${cst.blog_file}: ${err}. ${@FILE_LINE}')
	}

	defer {
		file.close()
	}

	emit_header(mut file, &b)!
}

fn parse_blog(lines []string) !Blog {
	mut topics := []TopicItem{}
	// mut locked := false

	if lines.len < 1 {
		return error('${cst.blog_file} is empty or incomplete. ${@FILE_LINE}')
	}

	name := util.parse_name_value('name=', lines[0]) or {
		return error('Unable to extract "name" from ${cst.blog_file}. ${@FILE_LINE}')
	}

	for i in 1 .. lines.len {
		t, dte, locked := util.parse_topic_values('topic', lines[i]) or {
			return error('util.parse_topic_values(...) returns nothing for line \'${lines[i]}\' in ${cst.blog_file} blog file. ${@FILE_LINE}')
		}
		topics << TopicItem{t, dte, locked}
	}
	return Blog{name, topics}
}

/**
 * This method generates topics's index page. It reads a fixed template, and ouput it as it it. When/If the
 * special tag is found, it inserts there, HTML code of links.
 */
pub fn (b &Blog) generate_topics_list_html() ! {
	// Open and load all post template file.
	mut t_lines := os.read_lines(cst.topics_list_template_file) or {
		return error('failed opening ${cst.topics_list_template_file} : ${err}. ${@FILE_LINE}\n [Tip: are you in the blog\'s root directory ?]')
	}

	// Copy Link model for later use. +1 to skip [LinkModel] tag
	link_model, lmt, em := util.extract_link_model(t_lines)!

	// Replace lines from [linkModel] to [EndModel] with Link tag: NOT OPTIMAL, IMPLIES MANY COPY
	t_lines.delete_many(lmt, em - lmt + 1)
	t_lines.insert(lmt, cst.list_links_tag)

	// Now create/overwrite output file
	mut index := os.open_file('${cst.topics_list_filename}', 'w+', cst.file_access) or {
		return error('opening ${cst.topics_list_filename} : ${err}. ${@FILE_LINE}\n [Tip: are you in the blog\'s root directory ?]')
	}

	defer {
		index.close()
	}

	mut dyn := util.DynVars.new()
	for l in t_lines {
		// replace potential DynVar in the line.
		dyn.add('@num', b.topics.len.str())
		s := dyn.substitute(l)!

		if s.contains(cst.list_links_tag) {
			// Emit all links
			for topic in b.topics {
				dir := util.obfuscate(topic.title)
				dyn.add('@url', '${dir}${os.path_separator}${cst.pushs_list_filename}')
				dyn.add('@title', topic.title)
				dyn.add('@date', util.to_blog_date(topic.date))

				// Emit full link model lines.
				for model_lines in link_model {
					f := dyn.substitute(model_lines)!
					index.writeln(f) or {
						return error('Unable to write ${cst.topics_list_filename}: ${err}. ${@FILE_LINE}')
					}
				}
			}
		} else {
			index.writeln(s) or {
				return error('Unable to write ${cst.topics_list_filename}: ${err}. ${@FILE_LINE}')
			}
		}
	}
}
