module commands

import term
import os
import constants as cst
import structures {Blog, Topic, Post}
import util

// Init structure, implementing Command interface.
struct Push implements Command {
	name    string
	desc    string
	help    string
	arg_min int
	arg_max int
	exec    fn (s []string) ! @[required]
}

// new builds a Init Command.
pub fn Push.new() Command {
	return Push{
		name:    'push'
		desc:    'Push a new article into topic (run from inside the topic directory).'
		help:    Push.help()
		arg_min: 1
		arg_max: 1
		exec:    push
	}
}

// help give a complete description of the command, including parameters.
fn Push.help() string {
	return '
Command: ${term.green('vssg')} ${term.yellow('push')} ${term.blue('path_to_text_file')}

The push command creates a new post in the current topic:

'
}

// push command feature are implemented here. The parameters number has been checked before call.
fn push(p []string) ! {
	post_file := p[0]

	// First, check post_file.
	if !os.exists('${post_file}') {
		return error('Error loading "${post_file}" : The file does not exist. ${@FILE_LINE}.')
	}


	mut topics := Topic.load()!
	id := topics.get_next_post_id()
	mut post := Post.load(post_file)!
	post.set_id(id)
	path := cst.push_dir_prefix + id.str()

	if os.exists('${path}') {
		return error('failed creating ${path} : The directory already exists. [${@FILE_LINE}]')
	}
	os.mkdir('./${path}', os.MkdirParams{0o755}) or { return error('mkdir ${path} fails: ${err}. [${@FILE_LINE}]') }
	println('Created push directory: ${term.blue(path)}')

	// Create a sub dir for pictures
	pic_dir := './${path}${os.path_separator}${cst.pushs_pic_dir}'
	os.mkdir(pic_dir, os.MkdirParams{0o755}) or { return error('mkdir ${pic_dir} fails: ${err}') }
	println('Created push images sub-directory :  ${term.blue(pic_dir)}')

}
