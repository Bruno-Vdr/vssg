module structures

import os
import io
import term
import time
import util
import constants as cst

// Structure that handle Post information, inside .topic file.
pub struct PostSummary {
pub:
	id    u64
	title string
	date  i64
	dir   string
}

pub struct Topic {
	title string // Topic title
pub:
	directory string // Dir. containing posts.
pub mut:
	posts []PostSummary
}

/**
 * Create a new empty topic, with no posts.
 */
pub fn Topic.new(title string) Topic {
	return Topic{title, util.obfuscate(title), []PostSummary{}}
}

/**
 * Load a topic file, removing comments and spaces at begining of lines.
 * Note: No parsing is done here, only strings loading.
 */
pub fn Topic.load() !Topic {
	mut ret := []string{} // []string is array type, []string{} declares an empty array.
	mut file := os.open(cst.topic_file) or {
		return error('Failed opening file ${cst.topic_file}: ${err}. [${@FILE_LINE}]\n[Hint: are you in the topics\'s directory ?]')
	}

	defer {
		file.close()
	}

	mut b_reader := io.new_buffered_reader(reader: file)
	for {
		mut s := b_reader.read_line() or { break }

		// Remove empty lines and comments # blabla
		s = s.trim_left(' ')
		if !s.starts_with('#') && s.len > 0 {
			ret << s
		}
	}
	return parse_topic_file(ret)!
}

fn parse_topic_file(lines []string) !Topic {
	mut posts := []PostSummary{}
	if lines.len == 0 {
		return error('${cst.topic_file} is empty. [${@FILE_LINE}]')
	}

	title := util.parse_name_value('topic=', lines[0]) or {
		return error('Unable to extract "title" from ${cst.topic_file}. [${@FILE_LINE}]')
	}

	directory := util.parse_name_value('directory=', lines[1]) or {
		return error('Unable to extract "directory" from ${cst.topic_file}. [${@FILE_LINE}]')
	}
	for i in 2 .. lines.len {
		id, t, date, dir := util.parse_push_values('push', lines[i]) or {
			return error('unable to parse "${lines[i]}". [${@FILE_LINE}]')
		}

		p := PostSummary{id, t, date, dir}
		posts << p
	}

	return Topic{title, directory, posts}
}

/**
 * Save Topic file containing posts relatives data.
 */
pub fn (t Topic) save(path string) ! {
	println('Updating ${cst.topic_file}  file in ./' + term.blue('${path}'))
	mut file := os.open_file('${path}${os.path_separator}${cst.topic_file}', 'w+', os.s_iwusr | os.s_irusr) or {
		return error('Unable to update $${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}

	defer {
		file.close()
	}
	date_time := time.now().str()
	file.writeln('#\n# Warning: do not edit this file ! It is dynamically generated by vssg.\n# Created on ${date_time} \n# This file contains Topic specific parameters (posts) for topic "${t.title}".\n#') or {
		return error('Unable to write ${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}
	file.writeln('topic="${t.title}"') or {
		return error('Unable to write ${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}
	file.writeln('directory="${t.directory}"') or {
		return error('Unable to write ${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}

	// Now list the defined posts
	for _, p in t.posts {
		file.writeln('push = [id:${p.id}][title:${p.title}][date:${p.date}][dir:.${os.path_separator}${cst.push_dir_prefix}${p.id}]') or {
			return error('Unable to write ${t.directory}${os.path_separator}${cst.topic_file}: ${err}, ${@FILE_LINE}')
		}
	}
}

pub fn (t Topic) get_next_post_id() u64 {
	// No entries at the moment. Next id is 0.
	if t.posts.len == 0 {
		return 0
	}

	mut next_id := u64(0)
	for p in t.posts {
		if p.id > next_id {
			next_id = p.id
		}
	}
	return next_id + 1
}

// This method generates posts index page. It reads a fixed template, and output it unchanged unless a dynamic
// variable is met or a special tag is found, it inserts there, HTML code of links.
pub fn (t Topic) generate_posts_list_html() ! {
	// Open post template file.
	mut t_lines := os.read_lines(cst.pushs_list_template_file) or {
		return error('Failed opening ${cst.pushs_list_template_file} : ${err}, ${@FILE_LINE}\n [Tip: are you in the Topic\'s directory ?]')
	}

	// Now extract [LinkModel]...[EndModel] section
	mut lmt := -1
	mut em := -1

	// Locate index of model tag start and stop.
	for i, l in t_lines {
		if l.contains(cst.link_model_tag) {
			lmt = i
		}
		if l.contains(cst.end_model) {
			em = i
		}
	}

	if lmt == -1 || em == -1 {
		return error('${cst.link_model_tag} or ${cst.end_model} tags not found in ${cst.pushs_list_template_file} template file. ${@FILE_LINE}')
	}

	if lmt >= em {
		return error('${cst.link_model_tag} or ${cst.end_model} order not respected in ${cst.pushs_list_template_file} template file. ${@FILE_LINE}')
	}

	// Copy Link model for later use. +1 to skip [LinkModel] tag
	link_model := t_lines[lmt + 1..em].clone()

	// Replace lines from [linkModel] to [EndModel] with Link tag: NOT OPTIMAL, IMPLIES MANY COPY
	t_lines.delete_many(lmt, em - lmt + 1)
	t_lines.insert(lmt, cst.list_links_tag)

	// Now create/overwrite output file
	mut index := os.open_file('${cst.pushs_list_filename}', 'w+', os.s_iwusr | os.s_irusr) or {
		return error('Error opening ${cst.pushs_list_filename} : ${err}, ${@FILE_LINE}\n [Tip: are you in the topics\'s directory ?]')
	}

	defer {
		index.close()
	}

	mut dyn := util.DynVars.new()
	for l in t_lines {
		// replace potential DynVar in the line.
		s := dyn.substitute(l)!

		if s.contains(cst.list_links_tag) {
			// Emit all links
			for post in t.posts {
				dir := cst.push_dir_prefix + post.id.str()
				dyn.add('@url', '${dir}${os.path_separator}${cst.push_filename}')
				dyn.add('@title', post.title)
				dyn.add('@date', util.to_blog_date(post.date))

				// Emit full link model lines.
				for model_lines in link_model {
					f := dyn.substitute(model_lines)!
					index.writeln(f) or {
						return error('Unable to write ${cst.pushs_list_filename}: ${err}, ${@FILE_LINE}')
					}
				}
			}
		} else {
			index.writeln(s) or {
				return error('Unable to write ${cst.pushs_list_filename}: ${err}, ${@FILE_LINE}')
			}
		}
	}
}
