module structures

import os
import term
import time
import util
import constants as cst

// Structure that handle Post information, inside .topic file.
pub struct PostSummary {
pub:
	id    u64
	title string
	date  i64
	dir   string
}

pub struct Topic {
pub:
	title     string // Topic title
	directory string // Dir. containing posts.
	locked    bool   // Is the topic locked ?
mut:
	posts map[u64]PostSummary
}

// Create a new empty topic, with no posts.
pub fn Topic.new(title string) Topic {
	return Topic{title, util.obfuscate(title), false, map[u64]PostSummary{}}
}

// build a new topic with existing posts.
pub fn Topic.build(title string, locked bool, posts map[u64]PostSummary) Topic {
	return Topic{title, util.obfuscate(title), locked, posts}
}

/**
 * Load a topic file, removing comments and spaces at beginning of lines.
 * Note: No parsing is done here, only strings loading.
 */
pub fn Topic.load() !Topic {
	if util.where_am_i() != .topic_dir {
		return error('Unable to load ${cst.topic_file}.\n[Hint: Are you in a Topic\'s directory ?]')
	}

	mut ret := util.load_transform_text_file(cst.topic_file, util.del_empty_and_comments)!
	return parse_topic_file(ret)!
}

fn parse_topic_file(lines []string) !Topic {
	mut posts := map[u64]PostSummary{}
	if lines.len == 0 {
		return error('${cst.topic_file} is empty. [${@FILE_LINE}]')
	}

	title := util.parse_name_value('topic=', lines[0]) or {
		return error('Unable to extract "title" from ${cst.topic_file}. [${@FILE_LINE}]')
	}

	directory := util.parse_name_value('directory=', lines[1]) or {
		return error('Unable to extract "directory" from ${cst.topic_file}. [${@FILE_LINE}]')
	}

	locked_str := util.parse_name_value('locked=', lines[2]) or {
		return error('Unable to extract "locked" from  "${lines[2]}" in ${cst.topic_file}. [${@FILE_LINE}]')
	}
	if locked_str !in ['true', 'false'] {
		return error('"locked" field is not true nor false in "${lines[2]}"')
	}

	locked := locked_str == 'true'

	for i in 3 .. lines.len {
		id, t, date, dir := util.parse_push_values('push', lines[i]) or {
			return error('unable to parse "${lines[i]}". [${@FILE_LINE}]')
		}

		p := PostSummary{id, t, date, dir}
		posts[p.id] = p
	}

	return Topic{title, directory, locked, posts}
}

/**
 * Save Topic file containing posts relatives data.
 */
pub fn (t Topic) save(path string) ! {
	println('Updating ${cst.topic_file}  file in ./' + term.blue('${path}'))
	mut file := os.open_file('${path}${os.path_separator}${cst.topic_file}', 'w+', cst.file_access) or {
		return error('Unable to update $${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}

	defer {
		file.close()
	}
	date_time := time.now().str()
	file.writeln('#\n# Warning: do not edit this file ! It is dynamically generated by vssg.\n# Created on ${date_time} \n# This file contains Topic specific parameters (posts) for topic "${t.title}".\n#') or {
		return error('Unable to write ${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}
	file.writeln('topic="${t.title}"') or {
		return error('Unable to write ${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}
	file.writeln('directory="${t.directory}"') or {
		return error('Unable to write ${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}
	file.writeln('locked="${t.locked}"') or {
		return error('Unable to write ${cst.topic_file}: ${err}, ${@FILE_LINE}')
	}

	// Now list the defined posts
	for _, p in t.posts {
		file.writeln('push = [id:${p.id}][title:${p.title}][date:${p.date}][dir:.${os.path_separator}${cst.push_dir_prefix}${p.id}]') or {
			return error('Unable to write ${t.directory}${os.path_separator}${cst.topic_file}: ${err}, ${@FILE_LINE}')
		}
	}
}

// get_posts_number return the number of post in the topic.
pub fn (t Topic) get_posts_number() int {
	return t.posts.len
}

// Return a COPY of the posts map
pub fn (t Topic) get_posts() map[u64]PostSummary {
	return t.posts.clone()
}

// Return PostSummary identified with id if any, none otherwise.
pub fn (t Topic) get_post(id u64) ?PostSummary {
	return if id in t.posts {
		t.posts[id]
	} else {
		none
	}
}

// Set/Add or Replace post based on its id. If id already exist, post is replace, else it's added.
pub fn (mut t Topic) set_post(ps PostSummary) {
	t.posts[ps.id] = ps
}

// delete a post from posts map, given the post id.
pub fn (mut t Topic) delete(id u64) ! {
	if id in t.posts {
		t.posts.delete(id)
	} else {
		return error('Non existing post with id=${id}.')
	}
}

pub fn (t Topic) get_next_post_id() u64 {
	// No entries at the moment. Next id is 0.
	if t.posts.len == 0 {
		return 0
	}

	mut next_id := u64(0)
	for _, v in t.posts {
		if v.id > next_id {
			next_id = v.id
		}
	}
	return next_id + 1
}

// get_last_post_summary return the last (highest) topic id, if any.
pub fn (t Topic) get_last_post_summary() ?PostSummary {
	if t.posts.len == 0 {
		return none
	} else {
		mut last_push := t.posts[0]
		for _, ps in t.posts {
			if ps.id > last_push.id {
				last_push = ps
			}
		}
		return last_push
	}
}

// This method generates pushs index page. It reads a fixed template, and output it unchanged unless a dynamic
// variable is met or a special tag is found, it inserts there, HTML code of links.
pub fn (t Topic) generate_pushes_list_html() ! {
	// Open post template file.
	mut t_lines := os.read_lines(cst.pushs_list_template_file) or {
		return error('Failed opening ${cst.pushs_list_template_file} : ${err}, ${@FILE_LINE}\n [Tip: are you in the Topic\'s directory ?]')
	}

	// Copy Link model for later use. +1 to skip [LinkModel] tag
	link_model, lmt, em := util.extract_link_model(t_lines)!

	// Replace lines from [linkModel] to [EndModel] with Link tag: NOT OPTIMAL, IMPLIES MANY COPY
	t_lines.delete_many(lmt, em - lmt + 1)
	t_lines.insert(lmt, cst.list_links_tag)

	// Now create/overwrite output file
	mut index := os.open_file('${cst.pushs_list_filename}', 'w+', cst.file_access) or {
		return error('Error opening ${cst.pushs_list_filename} : ${err}, ${@FILE_LINE}\n [Tip: are you in the topics\'s directory ?]')
	}

	defer {
		index.close()
	}

	mut dyn := util.DynVars.new()
	dyn.add('@topic', t.title)

	for l in t_lines {
		// replace potential DynVar in the line.
		dyn.add('@num', t.posts.len.str())
		s := dyn.substitute(l)!

		if s.contains(cst.list_links_tag) {
			// Emit all links
			for _, post in t.posts {
				dir := cst.push_dir_prefix + post.id.str()
				dyn.add('@url', '${dir}${os.path_separator}${cst.push_filename}')
				dyn.add('@title', post.title)
				dyn.add('@date', util.to_blog_date(post.date))
				dyn.add('@topic', t.title)

				// Emit full link model lines.
				for model_lines in link_model {
					f := dyn.substitute(model_lines)!
					index.writeln(f) or {
						return error('Unable to write ${cst.pushs_list_filename}: ${err}, ${@FILE_LINE}')
					}
				}
			}
		} else {
			index.writeln(s) or {
				return error('Unable to write ${cst.pushs_list_filename}: ${err}, ${@FILE_LINE}')
			}
		}
	}
}
