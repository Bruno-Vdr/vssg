module constants

pub const blog_file = '.blog'
pub const topic_file = '.topic'
