module structures

pub struct Blog {
}
