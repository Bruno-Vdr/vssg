module structures

import io
import os
import time
import term
import hash.fnv1a
import constants as cst
import util

/**
 * Blog contains arbitrary topic (subject/category/sub-section). This structure store the list of topics,
 * with title (shown) and creation date (time since epoq).
 */
pub struct Blog {
	name string
mut:
	topics []string
	date   []i64
}

// Static method to build empty Blog struct
pub fn Blog.new(name string) Blog {
	return Blog{name, []string{}, []i64{}}
}

// Static method that obfuscate a topic name
pub fn Blog.obfuscate(title string) string {
	return fnv1a.sum64_string(title).hex()
}

// Static method, loading blog file from current directory.
fn Blog.load() !Blog {
	mut ret := []string{} // []string is array type, []string{} declares an empty array.
	mut file := os.open(cst.blog_file) or {
		return error('opening file : ${err}\n[Hint: are you in the blog\'s root directory ?] ${@FILE_LINE}')
	}

	defer {
		file.close()
	}

	mut b_reader := io.new_buffered_reader(reader: file)
	for {
		mut s := b_reader.read_line() or { break }

		// Remove empty lines and comments # blabla
		s = s.trim_left(' ')
		if !s.starts_with('#') && s.len > 0 {
			ret << s
		}
	}

	return parse_blog(ret)
}

pub fn (mut b Blog) add_topic(topic string) {
	b.topics << topic
	b.date << time.ticks() / 1000 // Unix epoque in seconds !
}

pub fn (b Blog) get_topic(i int) ?(string, i64) {
	if i < b.topics.len {
		return b.topics[i], b.date[i]
	}
	return none
}

// Save the blog_file configuration.
pub fn (b Blog) save() ! {
	println('Updating ${cst.blog_file}  file in ' + term.blue('${b.name}'))
	mut file := os.open_file('${cst.blog_file}', 'w+', os.s_iwusr | os.s_irusr) or {
		return error('Unable to update ${cst.blog_file}: ${err}')
	}

	defer {
		file.close()
	}

	emit_header(mut file, b)!
	emit_topics(mut file, b)!
}

// emit_header write comments and  header only (no topics) int blog_file.
fn emit_header(mut file os.File, b &Blog) ! {
	date_time := time.now().str()
	file.writeln('#\n# Warning: do not edit this file ! It is dynamically generated by vssg.\n# Created on ${date_time} \n# This file contains blog specific parameters for "${b.name}".\n#') or {
		return error('Unable to write ${cst.blog_file}: ${err}')
	}

	file.writeln('name="${b.name}"') or {
		return error('Unable to write name in ${cst.blog_file}: ${err}')
	}
}

// emit_topics writes topics only into blog_file.
fn emit_topics(mut file os.File, b &Blog) ! {
	// Now list the defined topics
	for i, t in b.topics {
		file.writeln('topic="${t}" [${b.date[i]}] # In directory ./${b.name}/' + Blog.obfuscate(t)) or {
			return error('Unable to write ${cst.blog_file}: ${err}')
		}
	}
}

/**
 *  Create the initial blog file, containing only the name. At this time, no topics
 * have been added.
 * Note: This method is called in Init command, from outside the blog directory
 * so the configuration file is created with blog directory prepending. Other
 * commands are run from within the blog root's directory (to differentiate them) and
 * access to config_file don't need root's blog prefix.
 */
pub fn (b Blog) create() ! {
	println('Creating ${cst.blog_file}  file in ' + term.blue('${b.name}'))
	mut file := os.open_file('${b.name}${os.path_separator}${cst.blog_file}', 'w+', os.s_iwusr | os.s_irusr) or {
		return error('Unable to update ${b.name}${os.path_separator}${cst.blog_file}: ${err}. ${@FILE_LINE}')
	}

	defer {
		file.close()
	}

	emit_header(mut file, &b)!
}

fn parse_blog(lines []string) !Blog {
	mut topics := []string{}
	mut dates := []i64{}

	if lines.len < 1 {
		return error('Error: ${cst.blog_file} is empty or incomplete.')
	}

	name := util.parse_name_value('name=', lines[0]) or {
		return error('Unable to extract "name" from ${cst.blog_file}')
	}

	for i in 1 .. lines.len {
		t, dte := util.parse_topic_values('topic', lines[i]) or { return error('') }
		topics << t
		dates << dte
	}
	return Blog{name, topics, dates}
}

/**
 * This method generates topics's index page. It reads a fixed template, and ouput it as it it. When/If the
 * special tag is found, it inserts there, HTML code of links.
 */
fn (b &Blog) generate_topics_list_html() ! {
	// Open and load all post template file.
	mut t_lines := os.read_lines(cst.topics_list_template_file) or {
		return error('Error opening ${cst.topics_list_template_file} : ${err}\n [Tip: are you in the blog\'s root directory ?]')
	}

	// Now extract [LinkModel]...[EndModel] section
	mut lmt := -1
	mut em := -1

	// Locate index of model tag start and stop.
	for i, l in t_lines {
		if l.contains(cst.link_model_tag) {
			lmt = i
		}
		if l.contains(cst.end_model) {
			em = i
		}
	}

	if lmt == -1 || em == -1 {
		return error('${cst.link_model_tag} or ${cst.end_model} tags not found in ${cst.topics_list_template_file} template file.')
	}

	if lmt >= em {
		return error('${cst.link_model_tag} or ${cst.end_model} order not respected in ${cst.topics_list_template_file} template file.')
	}

	// Copy Link model for later use. +1 to skip [LinkModel] tag
	link_model := t_lines[lmt + 1..em].clone()

	// Replace lines from [linkModel] to [EndModel] with Link tag: NOT OPTIMAL, IMPLIES MANY COPY
	t_lines.delete_many(lmt, em - lmt + 1)
	t_lines.insert(lmt, cst.list_links_tag)

	// Now create/overwrite output file
	mut index := os.open_file('${cst.topics_list_filename}', 'w+', os.s_iwusr | os.s_irusr) or {
		return error('Error opening ${cst.topics_list_filename} : ${err}\n [Tip: are you in the blog\'s root directory ?]')
	}

	defer {
		index.close()
	}

	mut dyn := util.DynVars.new()
	for l in t_lines {
		// replace potential DynVar in the line.
		s := dyn.substitute(l)!

		if s.contains(cst.list_links_tag) {
			// Emit all links
			for i, topic in b.topics {
				dir := Blog.obfuscate(topic)
				dyn.add('@url', '${dir}${os.path_separator}${cst.posts_list_filename}')
				dyn.add('@title', b.topics[i])
				dyn.add('@date', util.to_blog_date(b.date[i]))

				// Emit full link model lines.
				for model_lines in link_model {
					f := dyn.substitute(model_lines)!
					index.writeln(f) or {
						return error('Unable to write ${cst.topics_list_filename}: ${err}')
					}
				}
			}
		} else {
			index.writeln(s) or {
				return error('Unable to write ${cst.topics_list_filename}: ${err}')
			}
		}
	}
}
